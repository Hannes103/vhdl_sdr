library ieee;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;

package iq_demodulator_pkg is
   
   type t_sfixed_array is array(natural range <>) of sfixed;
    
end package iq_demodulator_pkg;
